`include "transaction.sv"
`include "generator.sv"
`include "intf.sv"
`include "driver.sv"
`include "environment.sv"
`include "test.sv"
`include "design.v"
`include "assert_debounce.sv"
`include "testbench_top.sv"
