interface intf(input logic clk,reset);

logic sw;
logic db;

endinterface

